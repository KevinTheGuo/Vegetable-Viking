// nios_system.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module nios_system (
		input  wire        clk_clk,            //         clk.clk
		input  wire        reset_reset_n,      //       reset.reset_n
		output wire        sdram_clk_clk,      //   sdram_clk.clk
		output wire [12:0] sdram_wire_addr,    //  sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,      //            .ba
		output wire        sdram_wire_cas_n,   //            .cas_n
		output wire        sdram_wire_cke,     //            .cke
		output wire        sdram_wire_cs_n,    //            .cs_n
		inout  wire [31:0] sdram_wire_dq,      //            .dq
		output wire [3:0]  sdram_wire_dqm,     //            .dqm
		output wire        sdram_wire_ras_n,   //            .ras_n
		output wire        sdram_wire_we_n,    //            .we_n
		output wire [31:0] to_hw_port0_export, // to_hw_port0.export
		output wire [31:0] to_hw_port1_export, // to_hw_port1.export
		output wire [31:0] to_hw_port2_export, // to_hw_port2.export
		output wire [31:0] to_hw_port3_export, // to_hw_port3.export
		output wire [31:0] to_hw_port4_export, // to_hw_port4.export
		output wire [31:0] to_hw_port5_export, // to_hw_port5.export
		output wire [31:0] to_hw_port6_export, // to_hw_port6.export
		output wire [31:0] to_hw_port7_export, // to_hw_port7.export
		output wire [31:0] to_hw_port8_export, // to_hw_port8.export
		output wire [31:0] to_hw_port9_export, // to_hw_port9.export
		output wire [1:0]  to_hw_sig_export,   //   to_hw_sig.export
		input  wire [1:0]  to_sw_sig_export    //   to_sw_sig.export
	);

	wire         sdram_pll_c0_clk;                                            // sdram_pll:c0 -> [mm_interconnect_0:sdram_pll_c0_clk, rst_controller_002:clk, sdram:clk]
	wire  [31:0] nios2_qsys_0_data_master_readdata;                           // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire         nios2_qsys_0_data_master_debugaccess;                        // nios2_qsys_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire  [28:0] nios2_qsys_0_data_master_address;                            // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                         // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire         nios2_qsys_0_data_master_read;                               // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire         nios2_qsys_0_data_master_write;                              // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire  [31:0] nios2_qsys_0_data_master_writedata;                          // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire         nios2_qsys_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [28:0] nios2_qsys_0_instruction_master_address;                     // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                        // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;       // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;        // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_readdata;     // nios2_qsys_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_qsys_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_waitrequest;  // nios2_qsys_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_qsys_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_debugaccess -> nios2_qsys_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_address -> nios2_qsys_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_read -> nios2_qsys_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_byteenable -> nios2_qsys_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_write -> nios2_qsys_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_writedata -> nios2_qsys_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_readdata;              // sdram_pll:readdata -> mm_interconnect_0:sdram_pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_sdram_pll_pll_slave_address;               // mm_interconnect_0:sdram_pll_pll_slave_address -> sdram_pll:address
	wire         mm_interconnect_0_sdram_pll_pll_slave_read;                  // mm_interconnect_0:sdram_pll_pll_slave_read -> sdram_pll:read
	wire         mm_interconnect_0_sdram_pll_pll_slave_write;                 // mm_interconnect_0:sdram_pll_pll_slave_write -> sdram_pll:write
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_writedata;             // mm_interconnect_0:sdram_pll_pll_slave_writedata -> sdram_pll:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [15:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [2:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [1:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [15:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_sdram_s1_chipselect;                       // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                         // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                      // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                          // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                             // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                       // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                    // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                            // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                        // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_to_hw_port0_s1_chipselect;                 // mm_interconnect_0:to_hw_port0_s1_chipselect -> to_hw_port0:chipselect
	wire  [31:0] mm_interconnect_0_to_hw_port0_s1_readdata;                   // to_hw_port0:readdata -> mm_interconnect_0:to_hw_port0_s1_readdata
	wire   [1:0] mm_interconnect_0_to_hw_port0_s1_address;                    // mm_interconnect_0:to_hw_port0_s1_address -> to_hw_port0:address
	wire         mm_interconnect_0_to_hw_port0_s1_write;                      // mm_interconnect_0:to_hw_port0_s1_write -> to_hw_port0:write_n
	wire  [31:0] mm_interconnect_0_to_hw_port0_s1_writedata;                  // mm_interconnect_0:to_hw_port0_s1_writedata -> to_hw_port0:writedata
	wire         mm_interconnect_0_to_hw_port1_s1_chipselect;                 // mm_interconnect_0:to_hw_port1_s1_chipselect -> to_hw_port1:chipselect
	wire  [31:0] mm_interconnect_0_to_hw_port1_s1_readdata;                   // to_hw_port1:readdata -> mm_interconnect_0:to_hw_port1_s1_readdata
	wire   [1:0] mm_interconnect_0_to_hw_port1_s1_address;                    // mm_interconnect_0:to_hw_port1_s1_address -> to_hw_port1:address
	wire         mm_interconnect_0_to_hw_port1_s1_write;                      // mm_interconnect_0:to_hw_port1_s1_write -> to_hw_port1:write_n
	wire  [31:0] mm_interconnect_0_to_hw_port1_s1_writedata;                  // mm_interconnect_0:to_hw_port1_s1_writedata -> to_hw_port1:writedata
	wire         mm_interconnect_0_to_hw_port2_s1_chipselect;                 // mm_interconnect_0:to_hw_port2_s1_chipselect -> to_hw_port2:chipselect
	wire  [31:0] mm_interconnect_0_to_hw_port2_s1_readdata;                   // to_hw_port2:readdata -> mm_interconnect_0:to_hw_port2_s1_readdata
	wire   [1:0] mm_interconnect_0_to_hw_port2_s1_address;                    // mm_interconnect_0:to_hw_port2_s1_address -> to_hw_port2:address
	wire         mm_interconnect_0_to_hw_port2_s1_write;                      // mm_interconnect_0:to_hw_port2_s1_write -> to_hw_port2:write_n
	wire  [31:0] mm_interconnect_0_to_hw_port2_s1_writedata;                  // mm_interconnect_0:to_hw_port2_s1_writedata -> to_hw_port2:writedata
	wire         mm_interconnect_0_to_hw_port3_s1_chipselect;                 // mm_interconnect_0:to_hw_port3_s1_chipselect -> to_hw_port3:chipselect
	wire  [31:0] mm_interconnect_0_to_hw_port3_s1_readdata;                   // to_hw_port3:readdata -> mm_interconnect_0:to_hw_port3_s1_readdata
	wire   [1:0] mm_interconnect_0_to_hw_port3_s1_address;                    // mm_interconnect_0:to_hw_port3_s1_address -> to_hw_port3:address
	wire         mm_interconnect_0_to_hw_port3_s1_write;                      // mm_interconnect_0:to_hw_port3_s1_write -> to_hw_port3:write_n
	wire  [31:0] mm_interconnect_0_to_hw_port3_s1_writedata;                  // mm_interconnect_0:to_hw_port3_s1_writedata -> to_hw_port3:writedata
	wire         mm_interconnect_0_to_hw_port4_s1_chipselect;                 // mm_interconnect_0:to_hw_port4_s1_chipselect -> to_hw_port4:chipselect
	wire  [31:0] mm_interconnect_0_to_hw_port4_s1_readdata;                   // to_hw_port4:readdata -> mm_interconnect_0:to_hw_port4_s1_readdata
	wire   [1:0] mm_interconnect_0_to_hw_port4_s1_address;                    // mm_interconnect_0:to_hw_port4_s1_address -> to_hw_port4:address
	wire         mm_interconnect_0_to_hw_port4_s1_write;                      // mm_interconnect_0:to_hw_port4_s1_write -> to_hw_port4:write_n
	wire  [31:0] mm_interconnect_0_to_hw_port4_s1_writedata;                  // mm_interconnect_0:to_hw_port4_s1_writedata -> to_hw_port4:writedata
	wire         mm_interconnect_0_to_hw_port5_s1_chipselect;                 // mm_interconnect_0:to_hw_port5_s1_chipselect -> to_hw_port5:chipselect
	wire  [31:0] mm_interconnect_0_to_hw_port5_s1_readdata;                   // to_hw_port5:readdata -> mm_interconnect_0:to_hw_port5_s1_readdata
	wire   [1:0] mm_interconnect_0_to_hw_port5_s1_address;                    // mm_interconnect_0:to_hw_port5_s1_address -> to_hw_port5:address
	wire         mm_interconnect_0_to_hw_port5_s1_write;                      // mm_interconnect_0:to_hw_port5_s1_write -> to_hw_port5:write_n
	wire  [31:0] mm_interconnect_0_to_hw_port5_s1_writedata;                  // mm_interconnect_0:to_hw_port5_s1_writedata -> to_hw_port5:writedata
	wire         mm_interconnect_0_to_hw_port6_s1_chipselect;                 // mm_interconnect_0:to_hw_port6_s1_chipselect -> to_hw_port6:chipselect
	wire  [31:0] mm_interconnect_0_to_hw_port6_s1_readdata;                   // to_hw_port6:readdata -> mm_interconnect_0:to_hw_port6_s1_readdata
	wire   [1:0] mm_interconnect_0_to_hw_port6_s1_address;                    // mm_interconnect_0:to_hw_port6_s1_address -> to_hw_port6:address
	wire         mm_interconnect_0_to_hw_port6_s1_write;                      // mm_interconnect_0:to_hw_port6_s1_write -> to_hw_port6:write_n
	wire  [31:0] mm_interconnect_0_to_hw_port6_s1_writedata;                  // mm_interconnect_0:to_hw_port6_s1_writedata -> to_hw_port6:writedata
	wire         mm_interconnect_0_to_hw_port8_s1_chipselect;                 // mm_interconnect_0:to_hw_port8_s1_chipselect -> to_hw_port8:chipselect
	wire  [31:0] mm_interconnect_0_to_hw_port8_s1_readdata;                   // to_hw_port8:readdata -> mm_interconnect_0:to_hw_port8_s1_readdata
	wire   [1:0] mm_interconnect_0_to_hw_port8_s1_address;                    // mm_interconnect_0:to_hw_port8_s1_address -> to_hw_port8:address
	wire         mm_interconnect_0_to_hw_port8_s1_write;                      // mm_interconnect_0:to_hw_port8_s1_write -> to_hw_port8:write_n
	wire  [31:0] mm_interconnect_0_to_hw_port8_s1_writedata;                  // mm_interconnect_0:to_hw_port8_s1_writedata -> to_hw_port8:writedata
	wire         mm_interconnect_0_to_hw_port9_s1_chipselect;                 // mm_interconnect_0:to_hw_port9_s1_chipselect -> to_hw_port9:chipselect
	wire  [31:0] mm_interconnect_0_to_hw_port9_s1_readdata;                   // to_hw_port9:readdata -> mm_interconnect_0:to_hw_port9_s1_readdata
	wire   [1:0] mm_interconnect_0_to_hw_port9_s1_address;                    // mm_interconnect_0:to_hw_port9_s1_address -> to_hw_port9:address
	wire         mm_interconnect_0_to_hw_port9_s1_write;                      // mm_interconnect_0:to_hw_port9_s1_write -> to_hw_port9:write_n
	wire  [31:0] mm_interconnect_0_to_hw_port9_s1_writedata;                  // mm_interconnect_0:to_hw_port9_s1_writedata -> to_hw_port9:writedata
	wire         mm_interconnect_0_to_hw_sig_s1_chipselect;                   // mm_interconnect_0:to_hw_sig_s1_chipselect -> to_hw_sig:chipselect
	wire  [31:0] mm_interconnect_0_to_hw_sig_s1_readdata;                     // to_hw_sig:readdata -> mm_interconnect_0:to_hw_sig_s1_readdata
	wire   [1:0] mm_interconnect_0_to_hw_sig_s1_address;                      // mm_interconnect_0:to_hw_sig_s1_address -> to_hw_sig:address
	wire         mm_interconnect_0_to_hw_sig_s1_write;                        // mm_interconnect_0:to_hw_sig_s1_write -> to_hw_sig:write_n
	wire  [31:0] mm_interconnect_0_to_hw_sig_s1_writedata;                    // mm_interconnect_0:to_hw_sig_s1_writedata -> to_hw_sig:writedata
	wire         mm_interconnect_0_to_hw_port7_s1_chipselect;                 // mm_interconnect_0:to_hw_port7_s1_chipselect -> to_hw_port7:chipselect
	wire  [31:0] mm_interconnect_0_to_hw_port7_s1_readdata;                   // to_hw_port7:readdata -> mm_interconnect_0:to_hw_port7_s1_readdata
	wire   [1:0] mm_interconnect_0_to_hw_port7_s1_address;                    // mm_interconnect_0:to_hw_port7_s1_address -> to_hw_port7:address
	wire         mm_interconnect_0_to_hw_port7_s1_write;                      // mm_interconnect_0:to_hw_port7_s1_write -> to_hw_port7:write_n
	wire  [31:0] mm_interconnect_0_to_hw_port7_s1_writedata;                  // mm_interconnect_0:to_hw_port7_s1_writedata -> to_hw_port7:writedata
	wire  [31:0] mm_interconnect_0_to_sw_sig_s1_readdata;                     // to_sw_sig:readdata -> mm_interconnect_0:to_sw_sig_s1_readdata
	wire   [1:0] mm_interconnect_0_to_sw_sig_s1_address;                      // mm_interconnect_0:to_sw_sig_s1_address -> to_sw_sig:address
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_qsys_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_qsys_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_qsys_0_reset_reset_bridge_in_reset_reset, nios2_qsys_0:reset_n, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [nios2_qsys_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_qsys_0_debug_reset_request_reset;                      // nios2_qsys_0:debug_reset_request -> [rst_controller:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [mm_interconnect_0:sysid_qsys_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_translator_001:in_reset, sdram_pll:reset, sysid_qsys_0:reset_n, to_hw_port0:reset_n, to_hw_port1:reset_n, to_hw_port2:reset_n, to_hw_port3:reset_n, to_hw_port4:reset_n, to_hw_port5:reset_n, to_hw_port6:reset_n, to_hw_port7:reset_n, to_hw_port8:reset_n, to_hw_port9:reset_n, to_hw_sig:reset_n, to_sw_sig:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                      // rst_controller_001:reset_req -> [onchip_memory2_0:reset_req, rst_translator_001:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                          // rst_controller_002:reset_out -> [mm_interconnect_0:sdram_reset_reset_bridge_in_reset_reset, sdram:reset_n]

	nios_system_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	nios_system_nios2_qsys_0 nios2_qsys_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_qsys_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_qsys_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_qsys_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_qsys_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_qsys_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_qsys_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_qsys_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_qsys_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_qsys_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_qsys_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_qsys_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_qsys_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_qsys_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	nios_system_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)            //       .reset_req
	);

	nios_system_sdram sdram (
		.clk            (sdram_pll_c0_clk),                         //   clk.clk
		.reset_n        (~rst_controller_002_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	nios_system_sdram_pll sdram_pll (
		.clk       (clk_clk),                                         //       inclk_interface.clk
		.reset     (rst_controller_001_reset_out_reset),              // inclk_interface_reset.reset
		.read      (mm_interconnect_0_sdram_pll_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_sdram_pll_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_sdram_pll_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_sdram_pll_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_sdram_pll_pll_slave_writedata), //                      .writedata
		.c0        (sdram_pll_c0_clk),                                //                    c0.clk
		.c1        (sdram_clk_clk),                                   //                    c1.clk
		.areset    (),                                                //        areset_conduit.export
		.locked    (),                                                //        locked_conduit.export
		.phasedone ()                                                 //     phasedone_conduit.export
	);

	nios_system_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	nios_system_to_hw_port0 to_hw_port0 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_to_hw_port0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_to_hw_port0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_to_hw_port0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_to_hw_port0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_to_hw_port0_s1_readdata),   //                    .readdata
		.out_port   (to_hw_port0_export)                           // external_connection.export
	);

	nios_system_to_hw_port0 to_hw_port1 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_to_hw_port1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_to_hw_port1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_to_hw_port1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_to_hw_port1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_to_hw_port1_s1_readdata),   //                    .readdata
		.out_port   (to_hw_port1_export)                           // external_connection.export
	);

	nios_system_to_hw_port0 to_hw_port2 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_to_hw_port2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_to_hw_port2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_to_hw_port2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_to_hw_port2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_to_hw_port2_s1_readdata),   //                    .readdata
		.out_port   (to_hw_port2_export)                           // external_connection.export
	);

	nios_system_to_hw_port0 to_hw_port3 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_to_hw_port3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_to_hw_port3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_to_hw_port3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_to_hw_port3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_to_hw_port3_s1_readdata),   //                    .readdata
		.out_port   (to_hw_port3_export)                           // external_connection.export
	);

	nios_system_to_hw_port0 to_hw_port4 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_to_hw_port4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_to_hw_port4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_to_hw_port4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_to_hw_port4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_to_hw_port4_s1_readdata),   //                    .readdata
		.out_port   (to_hw_port4_export)                           // external_connection.export
	);

	nios_system_to_hw_port0 to_hw_port5 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_to_hw_port5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_to_hw_port5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_to_hw_port5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_to_hw_port5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_to_hw_port5_s1_readdata),   //                    .readdata
		.out_port   (to_hw_port5_export)                           // external_connection.export
	);

	nios_system_to_hw_port0 to_hw_port6 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_to_hw_port6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_to_hw_port6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_to_hw_port6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_to_hw_port6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_to_hw_port6_s1_readdata),   //                    .readdata
		.out_port   (to_hw_port6_export)                           // external_connection.export
	);

	nios_system_to_hw_port0 to_hw_port7 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_to_hw_port7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_to_hw_port7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_to_hw_port7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_to_hw_port7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_to_hw_port7_s1_readdata),   //                    .readdata
		.out_port   (to_hw_port7_export)                           // external_connection.export
	);

	nios_system_to_hw_port0 to_hw_port8 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_to_hw_port8_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_to_hw_port8_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_to_hw_port8_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_to_hw_port8_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_to_hw_port8_s1_readdata),   //                    .readdata
		.out_port   (to_hw_port8_export)                           // external_connection.export
	);

	nios_system_to_hw_port0 to_hw_port9 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_to_hw_port9_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_to_hw_port9_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_to_hw_port9_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_to_hw_port9_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_to_hw_port9_s1_readdata),   //                    .readdata
		.out_port   (to_hw_port9_export)                           // external_connection.export
	);

	nios_system_to_hw_sig to_hw_sig (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_to_hw_sig_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_to_hw_sig_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_to_hw_sig_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_to_hw_sig_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_to_hw_sig_s1_readdata),   //                    .readdata
		.out_port   (to_hw_sig_export)                           // external_connection.export
	);

	nios_system_to_sw_sig to_sw_sig (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_to_sw_sig_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_to_sw_sig_s1_readdata), //                    .readdata
		.in_port  (to_sw_sig_export)                         // external_connection.export
	);

	nios_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                     //                                clk_0_clk.clk
		.sdram_pll_c0_clk                               (sdram_pll_c0_clk),                                            //                             sdram_pll_c0.clk
		.nios2_qsys_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // nios2_qsys_0_reset_reset_bridge_in_reset.reset
		.sdram_reset_reset_bridge_in_reset_reset        (rst_controller_002_reset_out_reset),                          //        sdram_reset_reset_bridge_in_reset.reset
		.sysid_qsys_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // sysid_qsys_0_reset_reset_bridge_in_reset.reset
		.nios2_qsys_0_data_master_address               (nios2_qsys_0_data_master_address),                            //                 nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest           (nios2_qsys_0_data_master_waitrequest),                        //                                         .waitrequest
		.nios2_qsys_0_data_master_byteenable            (nios2_qsys_0_data_master_byteenable),                         //                                         .byteenable
		.nios2_qsys_0_data_master_read                  (nios2_qsys_0_data_master_read),                               //                                         .read
		.nios2_qsys_0_data_master_readdata              (nios2_qsys_0_data_master_readdata),                           //                                         .readdata
		.nios2_qsys_0_data_master_write                 (nios2_qsys_0_data_master_write),                              //                                         .write
		.nios2_qsys_0_data_master_writedata             (nios2_qsys_0_data_master_writedata),                          //                                         .writedata
		.nios2_qsys_0_data_master_debugaccess           (nios2_qsys_0_data_master_debugaccess),                        //                                         .debugaccess
		.nios2_qsys_0_instruction_master_address        (nios2_qsys_0_instruction_master_address),                     //          nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest    (nios2_qsys_0_instruction_master_waitrequest),                 //                                         .waitrequest
		.nios2_qsys_0_instruction_master_read           (nios2_qsys_0_instruction_master_read),                        //                                         .read
		.nios2_qsys_0_instruction_master_readdata       (nios2_qsys_0_instruction_master_readdata),                    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.nios2_qsys_0_debug_mem_slave_address           (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_address),      //             nios2_qsys_0_debug_mem_slave.address
		.nios2_qsys_0_debug_mem_slave_write             (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_write),        //                                         .write
		.nios2_qsys_0_debug_mem_slave_read              (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_read),         //                                         .read
		.nios2_qsys_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_readdata),     //                                         .readdata
		.nios2_qsys_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_writedata),    //                                         .writedata
		.nios2_qsys_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_byteenable),   //                                         .byteenable
		.nios2_qsys_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_waitrequest),  //                                         .waitrequest
		.nios2_qsys_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_debugaccess),  //                                         .debugaccess
		.onchip_memory2_0_s1_address                    (mm_interconnect_0_onchip_memory2_0_s1_address),               //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                         .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                         .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                         .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                         .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                         .clken
		.sdram_s1_address                               (mm_interconnect_0_sdram_s1_address),                          //                                 sdram_s1.address
		.sdram_s1_write                                 (mm_interconnect_0_sdram_s1_write),                            //                                         .write
		.sdram_s1_read                                  (mm_interconnect_0_sdram_s1_read),                             //                                         .read
		.sdram_s1_readdata                              (mm_interconnect_0_sdram_s1_readdata),                         //                                         .readdata
		.sdram_s1_writedata                             (mm_interconnect_0_sdram_s1_writedata),                        //                                         .writedata
		.sdram_s1_byteenable                            (mm_interconnect_0_sdram_s1_byteenable),                       //                                         .byteenable
		.sdram_s1_readdatavalid                         (mm_interconnect_0_sdram_s1_readdatavalid),                    //                                         .readdatavalid
		.sdram_s1_waitrequest                           (mm_interconnect_0_sdram_s1_waitrequest),                      //                                         .waitrequest
		.sdram_s1_chipselect                            (mm_interconnect_0_sdram_s1_chipselect),                       //                                         .chipselect
		.sdram_pll_pll_slave_address                    (mm_interconnect_0_sdram_pll_pll_slave_address),               //                      sdram_pll_pll_slave.address
		.sdram_pll_pll_slave_write                      (mm_interconnect_0_sdram_pll_pll_slave_write),                 //                                         .write
		.sdram_pll_pll_slave_read                       (mm_interconnect_0_sdram_pll_pll_slave_read),                  //                                         .read
		.sdram_pll_pll_slave_readdata                   (mm_interconnect_0_sdram_pll_pll_slave_readdata),              //                                         .readdata
		.sdram_pll_pll_slave_writedata                  (mm_interconnect_0_sdram_pll_pll_slave_writedata),             //                                         .writedata
		.sysid_qsys_0_control_slave_address             (mm_interconnect_0_sysid_qsys_0_control_slave_address),        //               sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata            (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),       //                                         .readdata
		.to_hw_port0_s1_address                         (mm_interconnect_0_to_hw_port0_s1_address),                    //                           to_hw_port0_s1.address
		.to_hw_port0_s1_write                           (mm_interconnect_0_to_hw_port0_s1_write),                      //                                         .write
		.to_hw_port0_s1_readdata                        (mm_interconnect_0_to_hw_port0_s1_readdata),                   //                                         .readdata
		.to_hw_port0_s1_writedata                       (mm_interconnect_0_to_hw_port0_s1_writedata),                  //                                         .writedata
		.to_hw_port0_s1_chipselect                      (mm_interconnect_0_to_hw_port0_s1_chipselect),                 //                                         .chipselect
		.to_hw_port1_s1_address                         (mm_interconnect_0_to_hw_port1_s1_address),                    //                           to_hw_port1_s1.address
		.to_hw_port1_s1_write                           (mm_interconnect_0_to_hw_port1_s1_write),                      //                                         .write
		.to_hw_port1_s1_readdata                        (mm_interconnect_0_to_hw_port1_s1_readdata),                   //                                         .readdata
		.to_hw_port1_s1_writedata                       (mm_interconnect_0_to_hw_port1_s1_writedata),                  //                                         .writedata
		.to_hw_port1_s1_chipselect                      (mm_interconnect_0_to_hw_port1_s1_chipselect),                 //                                         .chipselect
		.to_hw_port2_s1_address                         (mm_interconnect_0_to_hw_port2_s1_address),                    //                           to_hw_port2_s1.address
		.to_hw_port2_s1_write                           (mm_interconnect_0_to_hw_port2_s1_write),                      //                                         .write
		.to_hw_port2_s1_readdata                        (mm_interconnect_0_to_hw_port2_s1_readdata),                   //                                         .readdata
		.to_hw_port2_s1_writedata                       (mm_interconnect_0_to_hw_port2_s1_writedata),                  //                                         .writedata
		.to_hw_port2_s1_chipselect                      (mm_interconnect_0_to_hw_port2_s1_chipselect),                 //                                         .chipselect
		.to_hw_port3_s1_address                         (mm_interconnect_0_to_hw_port3_s1_address),                    //                           to_hw_port3_s1.address
		.to_hw_port3_s1_write                           (mm_interconnect_0_to_hw_port3_s1_write),                      //                                         .write
		.to_hw_port3_s1_readdata                        (mm_interconnect_0_to_hw_port3_s1_readdata),                   //                                         .readdata
		.to_hw_port3_s1_writedata                       (mm_interconnect_0_to_hw_port3_s1_writedata),                  //                                         .writedata
		.to_hw_port3_s1_chipselect                      (mm_interconnect_0_to_hw_port3_s1_chipselect),                 //                                         .chipselect
		.to_hw_port4_s1_address                         (mm_interconnect_0_to_hw_port4_s1_address),                    //                           to_hw_port4_s1.address
		.to_hw_port4_s1_write                           (mm_interconnect_0_to_hw_port4_s1_write),                      //                                         .write
		.to_hw_port4_s1_readdata                        (mm_interconnect_0_to_hw_port4_s1_readdata),                   //                                         .readdata
		.to_hw_port4_s1_writedata                       (mm_interconnect_0_to_hw_port4_s1_writedata),                  //                                         .writedata
		.to_hw_port4_s1_chipselect                      (mm_interconnect_0_to_hw_port4_s1_chipselect),                 //                                         .chipselect
		.to_hw_port5_s1_address                         (mm_interconnect_0_to_hw_port5_s1_address),                    //                           to_hw_port5_s1.address
		.to_hw_port5_s1_write                           (mm_interconnect_0_to_hw_port5_s1_write),                      //                                         .write
		.to_hw_port5_s1_readdata                        (mm_interconnect_0_to_hw_port5_s1_readdata),                   //                                         .readdata
		.to_hw_port5_s1_writedata                       (mm_interconnect_0_to_hw_port5_s1_writedata),                  //                                         .writedata
		.to_hw_port5_s1_chipselect                      (mm_interconnect_0_to_hw_port5_s1_chipselect),                 //                                         .chipselect
		.to_hw_port6_s1_address                         (mm_interconnect_0_to_hw_port6_s1_address),                    //                           to_hw_port6_s1.address
		.to_hw_port6_s1_write                           (mm_interconnect_0_to_hw_port6_s1_write),                      //                                         .write
		.to_hw_port6_s1_readdata                        (mm_interconnect_0_to_hw_port6_s1_readdata),                   //                                         .readdata
		.to_hw_port6_s1_writedata                       (mm_interconnect_0_to_hw_port6_s1_writedata),                  //                                         .writedata
		.to_hw_port6_s1_chipselect                      (mm_interconnect_0_to_hw_port6_s1_chipselect),                 //                                         .chipselect
		.to_hw_port7_s1_address                         (mm_interconnect_0_to_hw_port7_s1_address),                    //                           to_hw_port7_s1.address
		.to_hw_port7_s1_write                           (mm_interconnect_0_to_hw_port7_s1_write),                      //                                         .write
		.to_hw_port7_s1_readdata                        (mm_interconnect_0_to_hw_port7_s1_readdata),                   //                                         .readdata
		.to_hw_port7_s1_writedata                       (mm_interconnect_0_to_hw_port7_s1_writedata),                  //                                         .writedata
		.to_hw_port7_s1_chipselect                      (mm_interconnect_0_to_hw_port7_s1_chipselect),                 //                                         .chipselect
		.to_hw_port8_s1_address                         (mm_interconnect_0_to_hw_port8_s1_address),                    //                           to_hw_port8_s1.address
		.to_hw_port8_s1_write                           (mm_interconnect_0_to_hw_port8_s1_write),                      //                                         .write
		.to_hw_port8_s1_readdata                        (mm_interconnect_0_to_hw_port8_s1_readdata),                   //                                         .readdata
		.to_hw_port8_s1_writedata                       (mm_interconnect_0_to_hw_port8_s1_writedata),                  //                                         .writedata
		.to_hw_port8_s1_chipselect                      (mm_interconnect_0_to_hw_port8_s1_chipselect),                 //                                         .chipselect
		.to_hw_port9_s1_address                         (mm_interconnect_0_to_hw_port9_s1_address),                    //                           to_hw_port9_s1.address
		.to_hw_port9_s1_write                           (mm_interconnect_0_to_hw_port9_s1_write),                      //                                         .write
		.to_hw_port9_s1_readdata                        (mm_interconnect_0_to_hw_port9_s1_readdata),                   //                                         .readdata
		.to_hw_port9_s1_writedata                       (mm_interconnect_0_to_hw_port9_s1_writedata),                  //                                         .writedata
		.to_hw_port9_s1_chipselect                      (mm_interconnect_0_to_hw_port9_s1_chipselect),                 //                                         .chipselect
		.to_hw_sig_s1_address                           (mm_interconnect_0_to_hw_sig_s1_address),                      //                             to_hw_sig_s1.address
		.to_hw_sig_s1_write                             (mm_interconnect_0_to_hw_sig_s1_write),                        //                                         .write
		.to_hw_sig_s1_readdata                          (mm_interconnect_0_to_hw_sig_s1_readdata),                     //                                         .readdata
		.to_hw_sig_s1_writedata                         (mm_interconnect_0_to_hw_sig_s1_writedata),                    //                                         .writedata
		.to_hw_sig_s1_chipselect                        (mm_interconnect_0_to_hw_sig_s1_chipselect),                   //                                         .chipselect
		.to_sw_sig_s1_address                           (mm_interconnect_0_to_sw_sig_s1_address),                      //                             to_sw_sig_s1.address
		.to_sw_sig_s1_readdata                          (mm_interconnect_0_to_sw_sig_s1_readdata)                      //                                         .readdata
	);

	nios_system_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_qsys_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_qsys_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_qsys_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (sdram_pll_c0_clk),                       //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
